module main;
initial $interact;
endmodule
